module cpu(input instruction,
                 clk,
                 rst,
           output [31:0] pc);

    reg [31:0] pc;

    reg [

endmodule
